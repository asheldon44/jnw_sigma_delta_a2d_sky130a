*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/JNW_SIGMA_DELTA_A2D_lpe.spi
#else
.include ../../../work/xsch/JNW_SIGMA_DELTA_A2D.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-4

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p
.param vdd = 1.8
.param AVDD = 1.8
.param per = 1/16e6

.model mysw SW vt{vdd/2} ron=10k roff=1gig"

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
V_ground  VSS  0     dc 0
V_sup  VDD_1V8  VSS  dc {AVDD}
V_IN IN VSS dc {vdd/2} sin({vdd/2} {vdd/4} 100k 1n 0 0)

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------
.save xdut.q xdut.qn xdut.res xdut.resb xdut.vcmp xdut.p1 xdut.p2 xdut.vo1 xdut.vo2

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

op

tran 0.25n 100u
write
quit

.endc

.end
